`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/01/12 20:52:46
// Design Name: 
// Module Name: getaddr
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module getaddr(aclk,x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,
addra0,addra1,addra2,addra3,addra4,addra5,addra6,addra7,addra8,addra9,
addrb0,addrb1,addrb2,addrb3,addrb4,addrb5,addrb6,addrb7,addrb8,addrb9);
input aclk;
input [15:0] x0,x1,x2,x3,x4,x5,x6,x7,x8,x9;
output[5:0] addra0,addra1,addra2,addra3,addra4,addra5,addra6,addra7,addra8,addra9;
output[5:0] addrb0,addrb1,addrb2,addrb3,addrb4,addrb5,addrb6,addrb7,addrb8,addrb9;
reg [5:0] addra0,addra1,addra2,addra3,addra4,addra5,addra6,addra7,addra8,addra9;
reg [5:0] addrb0,addrb1,addrb2,addrb3,addrb4,addrb5,addrb6,addrb7,addrb8,addrb9;
always @(posedge aclk)
begin
if(x0[15:15]==1) //minus
        begin
        if((x0[14:0]<=15'b100100010000000)&&(x0[14:0]>15'b100100000000000)) //18560   18432
            begin
                addra0=6'b000000;
                addrb0=6'b000001;
            end
        else if((x0[14:0]<=15'b100100000000000)&&(x0[14:0]>15'b100011100000000)) //18432  18176
            begin
                addra0=6'b000010;
                addrb0=6'b000011;
            end
        else if((x0[14:0]<=15'b100011100000000)&&(x0[14:0]>15'b100011000000000))//18176  17920
            begin
                addra0=6'b000100;
                addrb0=6'b000101;
            end
        else if((x0[14:0]<=15'b100011000000000)&&(x0[14:0]>15'b100010100000000))
            begin
                addra0=6'b000110;
                addrb0=6'b000111;
            end
        else if((x0[14:0]<=15'b100010100000000)&&(x0[14:0]>15'b100010000000000))
            begin
                addra0=6'b001000;
                addrb0=6'b001001;
            end
        else if((x0[14:0]<=15'b100010000000000)&&(x0[14:0]>15'b100001000000000))
            begin
                addra0=6'b001010;
                addrb0=6'b001011;
            end
        else if((x0[14:0]<=15'b100001000000000)&&(x0[14:0]>15'b100000000000000))
            begin
                addra0=6'b001100;
                addrb0=6'b001101;
            end
        else if((x0[14:0]<=15'b100000000000000)&&(x0[14:0]>15'b011110000000000))
            begin
                addra0=6'b001110;
                addrb0=6'b001111;
            end
        else if((x0[14:0]<=15'b011110000000000)&&(x0[14:0]>15'b000000000000000))
            begin
                addra0=6'b010000;
                addrb0=6'b010001;
            end
            end
else
     begin
        if((x0[14:0]<=15'b011110000000000)&&(x0[14:0]>15'b000000000000000))
            begin
                addra0=6'b010010;
                addrb0=6'b010011;
            end
        else if((x0[14:0]<=15'b100000000000000)&&(x0>15'b011110000000000))
            begin
                addra0=6'b010100;
                addrb0=6'b010101;
            end
        else if((x0[14:0]<=15'b100001000000000)&&(x0>15'b100000000000000))
            begin
                addra0=6'b010110;
                addrb0=6'b010111;
            end
        else if((x0[14:0]<=15'b100010000000000)&&(x0[14:0]>15'b100001000000000))
            begin
                addra0=6'b011000;
                addrb0=6'b011001;
            end
        else if((x0[14:0]<=15'b100010100000000)&&(x0[14:0]>15'b100010000000000))
            begin
                addra0=6'b011010;
                addrb0=6'b011011;
            end
        else if((x0[14:0]<=15'b100011000000000)&&(x0[14:0]>15'b100010100000000))
            begin
                addra0=6'b011100;
                addrb0=6'b011101;
            end
        else if((x0[14:0]<=15'b100011100000000)&&(x0[14:0]>15'b100011000000000))
            begin
                addra0=6'b011110;
                addrb0=6'b011111;
            end
        else if((x0[14:0]<=15'b100100000000000)&&(x0[14:0]>15'b100011100000000))
            begin
                addra0=6'b100000;
                addrb0=6'b100001;
            end
        else if((x0[14:0]<=15'b100100010000000)&&(x0[14:0]>15'b100100000000000))
            begin
                addra0=6'b100010;
                addrb0=6'b100011;
            end
        else if((x0[14:0]<=15'b100100100000000)&&(x0[14:0]>15'b100100010000000))
            begin
                addra0=6'b100100;
                addrb0=6'b100101;
            end
    end
    end
always @(posedge aclk)
    begin
    if(x1[15:15]==1)
            begin
            if((x1[14:0]<=15'b100100010000000)&&(x1[14:0]>15'b100100000000000)) 
                begin
                    addra1=6'b000000;
                    addrb1=6'b000001;
                end
            else if((x1[14:0]<=15'b100100000000000)&&(x1[14:0]>15'b100011100000000))
                begin
                    addra1=6'b000010;
                    addrb1=6'b000011;
                end
            else if((x1[14:0]<=15'b100011100000000)&&(x1[14:0]>15'b100011000000000))
                begin
                    addra1=6'b000100;
                    addrb1=6'b000101;
                end
            else if((x1[14:0]<=15'b100011000000000)&&(x1[14:0]>15'b100010100000000))
                begin
                    addra1=6'b000110;
                    addrb1=6'b000111;
                end
            else if((x1[14:0]<=15'b100010100000000)&&(x1[14:0]>15'b100010000000000))
                begin
                    addra1=6'b001000;
                    addrb1=6'b001001;
                end
            else if((x1[14:0]<=15'b100010000000000)&&(x1[14:0]>15'b100001000000000))
                begin
                    addra1=6'b001010;
                    addrb1=6'b001011;
                end
            else if((x1[14:0]<=15'b100001000000000)&&(x1[14:0]>15'b100000000000000))
                begin
                    addra1=6'b001100;
                    addrb1=6'b001101;
                end
            else if((x1[14:0]<=15'b100000000000000)&&(x1[14:0]>15'b011110000000000))
                begin
                    addra1=6'b001110;
                    addrb1=6'b001111;
                end
            else if((x1[14:0]<=15'b011110000000000)&&(x1[14:0]>15'b000000000000000))
                begin
                    addra1=6'b010000;
                    addrb1=6'b010001;
                end
                end
    else
         begin
            if((x1[14:0]<=15'b011110000000000)&&(x1[14:0]>15'b000000000000000))
                begin
                    addra1=6'b010010;
                    addrb1=6'b010011;
                end
            else if((x1[14:0]<=15'b100000000000000)&&(x1>15'b011110000000000))
                begin
                    addra1=6'b010100;
                    addrb1=6'b010101;
                end
            else if((x1[14:0]<=15'b100001000000000)&&(x1>15'b100000000000000))
                begin
                    addra1=6'b010110;
                    addrb1=6'b010111;
                end
            else if((x1[14:0]<=15'b100010000000000)&&(x1[14:0]>15'b100001000000000))
                begin
                    addra1=6'b011000;
                    addrb1=6'b011001;
                end
            else if((x1[14:0]<=15'b100010100000000)&&(x1[14:0]>15'b100010000000000))
                begin
                    addra1=6'b011010;
                    addrb1=6'b011011;
                end
            else if((x1[14:0]<=15'b100011000000000)&&(x1[14:0]>15'b100010100000000))
                begin
                    addra1=6'b011100;
                    addrb1=6'b011101;
                end
            else if((x1[14:0]<=15'b100011100000000)&&(x1[14:0]>15'b100011000000000))
                begin
                    addra1=6'b011110;
                    addrb1=6'b011111;
                end
            else if((x1[14:0]<=15'b100100000000000)&&(x1[14:0]>15'b100011100000000))
                begin
                    addra1=6'b100000;
                    addrb1=6'b100001;
                end
            else if((x1[14:0]<=15'b100100010000000)&&(x1[14:0]>15'b100100000000000))
                begin
                    addra1=6'b100010;
                    addrb1=6'b100011;
                end
            else if((x1[14:0]<=15'b100100100000000)&&(x1[14:0]>15'b100100010000000))
                begin
                    addra1=6'b100100;
                    addrb1=6'b100101;
                end
        end
        end
    always @(posedge aclk)
    begin
    if(x2[15:15]==1)
            begin
            if((x2[14:0]<=15'b100100010000000)&&(x2[14:0]>15'b100100000000000)) 
                begin
                    addra2=6'b000000;
                    addrb2=6'b000001;
                end
            else if((x2[14:0]<=15'b100100000000000)&&(x2[14:0]>15'b100011100000000))
                begin
                    addra2=6'b000010;
                    addrb2=6'b000011;
                end
            else if((x2[14:0]<=15'b100011100000000)&&(x2[14:0]>15'b100011000000000))
                begin
                    addra2=6'b000100;
                    addrb2=6'b000101;
                end
            else if((x2[14:0]<=15'b100011000000000)&&(x2[14:0]>15'b100010100000000))
                begin
                    addra2=6'b000110;
                    addrb2=6'b000111;
                end
            else if((x2[14:0]<=15'b100010100000000)&&(x2[14:0]>15'b100010000000000))
                begin
                    addra2=6'b001000;
                    addrb2=6'b001001;
                end
            else if((x2[14:0]<=15'b100010000000000)&&(x2[14:0]>15'b100001000000000))
                begin
                    addra2=6'b001010;
                    addrb2=6'b001011;
                end
            else if((x2[14:0]<=15'b100001000000000)&&(x2[14:0]>15'b100000000000000))
                begin
                    addra2=6'b001100;
                    addrb2=6'b001101;
                end
            else if((x2[14:0]<=15'b100000000000000)&&(x2[14:0]>15'b011110000000000))
                begin
                    addra2=6'b001110;
                    addrb2=6'b001111;
                end
            else if((x2[14:0]<=15'b011110000000000)&&(x2[14:0]>15'b000000000000000))
                begin
                    addra2=6'b010000;
                    addrb2=6'b010001;
                end
                end
    else
         begin
            if((x2[14:0]<=15'b011110000000000)&&(x2[14:0]>15'b000000000000000))
                begin
                    addra2=6'b010010;
                    addrb2=6'b010011;
                end
            else if((x2[14:0]<=15'b100000000000000)&&(x2>15'b011110000000000))
                begin
                    addra2=6'b010100;
                    addrb2=6'b010101;
                end
            else if((x2[14:0]<=15'b100001000000000)&&(x2>15'b100000000000000))
                begin
                    addra2=6'b010110;
                    addrb2=6'b010111;
                end
            else if((x2[14:0]<=15'b100010000000000)&&(x2[14:0]>15'b100001000000000))
                begin
                    addra2=6'b011000;
                    addrb2=6'b011001;
                end
            else if((x2[14:0]<=15'b100010100000000)&&(x2[14:0]>15'b100010000000000))
                begin
                    addra2=6'b011010;
                    addrb2=6'b011011;
                end
            else if((x2[14:0]<=15'b100011000000000)&&(x2[14:0]>15'b100010100000000))
                begin
                    addra2=6'b011100;
                    addrb2=6'b011101;
                end
            else if((x2[14:0]<=15'b100011100000000)&&(x2[14:0]>15'b100011000000000))
                begin
                    addra2=6'b011110;
                    addrb2=6'b011111;
                end
            else if((x2[14:0]<=15'b100100000000000)&&(x2[14:0]>15'b100011100000000))
                begin
                    addra2=6'b100000;
                    addrb2=6'b100001;
                end
            else if((x2[14:0]<=15'b100100010000000)&&(x2[14:0]>15'b100100000000000))
                begin
                    addra2=6'b100010;
                    addrb2=6'b100011;
                end
            else if((x2[14:0]<=15'b100100100000000)&&(x2[14:0]>15'b100100010000000))
                begin
                    addra2=6'b100100;
                    addrb2=6'b100101;
                end
        end
        end
        always @(posedge aclk)
    begin
    if(x3[15:15]==1)
            begin
            if((x3[14:0]<=15'b100100010000000)&&(x3[14:0]>15'b100100000000000)) 
                begin
                    addra3=6'b000000;
                    addrb3=6'b000001;
                end
            else if((x3[14:0]<=15'b100100000000000)&&(x3[14:0]>15'b100011100000000))
                begin
                    addra3=6'b000010;
                    addrb3=6'b000011;
                end
            else if((x3[14:0]<=15'b100011100000000)&&(x3[14:0]>15'b100011000000000))
                begin
                    addra3=6'b000100;
                    addrb3=6'b000101;
                end
            else if((x3[14:0]<=15'b100011000000000)&&(x3[14:0]>15'b100010100000000))
                begin
                    addra3=6'b000110;
                    addrb3=6'b000111;
                end
            else if((x3[14:0]<=15'b100010100000000)&&(x3[14:0]>15'b100010000000000))
                begin
                    addra3=6'b001000;
                    addrb3=6'b001001;
                end
            else if((x3[14:0]<=15'b100010000000000)&&(x3[14:0]>15'b100001000000000))
                begin
                    addra3=6'b001010;
                    addrb3=6'b001011;
                end
            else if((x3[14:0]<=15'b100001000000000)&&(x3[14:0]>15'b100000000000000))
                begin
                    addra3=6'b001100;
                    addrb3=6'b001101;
                end
            else if((x3[14:0]<=15'b100000000000000)&&(x3[14:0]>15'b011110000000000))
                begin
                    addra3=6'b001110;
                    addrb3=6'b001111;
                end
            else if((x3[14:0]<=15'b011110000000000)&&(x3[14:0]>15'b000000000000000))
                begin
                    addra3=6'b010000;
                    addrb3=6'b010001;
                end
                end
    else
         begin
            if((x3[14:0]<=15'b011110000000000)&&(x3[14:0]>15'b000000000000000))
                begin
                    addra3=6'b010010;
                    addrb3=6'b010011;
                end
            else if((x3[14:0]<=15'b100000000000000)&&(x3>15'b011110000000000))
                begin
                    addra3=6'b010100;
                    addrb3=6'b010101;
                end
            else if((x3[14:0]<=15'b100001000000000)&&(x3>15'b100000000000000))
                begin
                    addra3=6'b010110;
                    addrb3=6'b010111;
                end
            else if((x3[14:0]<=15'b100010000000000)&&(x3[14:0]>15'b100001000000000))
                begin
                    addra3=6'b011000;
                    addrb3=6'b011001;
                end
            else if((x3[14:0]<=15'b100010100000000)&&(x3[14:0]>15'b100010000000000))
                begin
                    addra3=6'b011010;
                    addrb3=6'b011011;
                end
            else if((x3[14:0]<=15'b100011000000000)&&(x3[14:0]>15'b100010100000000))
                begin
                    addra3=6'b011100;
                    addrb3=6'b011101;
                end
            else if((x3[14:0]<=15'b100011100000000)&&(x3[14:0]>15'b100011000000000))
                begin
                    addra3=6'b011110;
                    addrb3=6'b011111;
                end
            else if((x3[14:0]<=15'b100100000000000)&&(x3[14:0]>15'b100011100000000))
                begin
                    addra3=6'b100000;
                    addrb3=6'b100001;
                end
            else if((x3[14:0]<=15'b100100010000000)&&(x3[14:0]>15'b100100000000000))
                begin
                    addra3=6'b100010;
                    addrb3=6'b100011;
                end
            else if((x3[14:0]<=15'b100100100000000)&&(x3[14:0]>15'b100100010000000))
                begin
                    addra3=6'b100100;
                    addrb3=6'b100101;
                end
        end
        end
        always @(posedge aclk)
    begin
    if(x4[15:15]==1)
            begin
            if((x4[14:0]<=15'b100100010000000)&&(x4[14:0]>15'b100100000000000)) 
                begin
                    addra4=6'b000000;
                    addrb4=6'b000001;
                end
            else if((x4[14:0]<=15'b100100000000000)&&(x4[14:0]>15'b100011100000000))
                begin
                    addra4=6'b000010;
                    addrb4=6'b000011;
                end
            else if((x4[14:0]<=15'b100011100000000)&&(x4[14:0]>15'b100011000000000))
                begin
                    addra4=6'b000100;
                    addrb4=6'b000101;
                end
            else if((x4[14:0]<=15'b100011000000000)&&(x4[14:0]>15'b100010100000000))
                begin
                    addra4=6'b000110;
                    addrb4=6'b000111;
                end
            else if((x4[14:0]<=15'b100010100000000)&&(x4[14:0]>15'b100010000000000))
                begin
                    addra4=6'b001000;
                    addrb4=6'b001001;
                end
            else if((x4[14:0]<=15'b100010000000000)&&(x4[14:0]>15'b100001000000000))
                begin
                    addra4=6'b001010;
                    addrb4=6'b001011;
                end
            else if((x4[14:0]<=15'b100001000000000)&&(x4[14:0]>15'b100000000000000))
                begin
                    addra4=6'b001100;
                    addrb4=6'b001101;
                end
            else if((x4[14:0]<=15'b100000000000000)&&(x4[14:0]>15'b011110000000000))
                begin
                    addra4=6'b001110;
                    addrb4=6'b001111;
                end
            else if((x4[14:0]<=15'b011110000000000)&&(x4[14:0]>15'b000000000000000))
                begin
                    addra4=6'b010000;
                    addrb4=6'b010001;
                end
                end
    else
         begin
            if((x4[14:0]<=15'b011110000000000)&&(x4[14:0]>15'b000000000000000))
                begin
                    addra4=6'b010010;
                    addrb4=6'b010011;
                end
            else if((x4[14:0]<=15'b100000000000000)&&(x4>15'b011110000000000))
                begin
                    addra4=6'b010100;
                    addrb4=6'b010101;
                end
            else if((x4[14:0]<=15'b100001000000000)&&(x4>15'b100000000000000))
                begin
                    addra4=6'b010110;
                    addrb4=6'b010111;
                end
            else if((x4[14:0]<=15'b100010000000000)&&(x4[14:0]>15'b100001000000000))
                begin
                    addra4=6'b011000;
                    addrb4=6'b011001;
                end
            else if((x4[14:0]<=15'b100010100000000)&&(x4[14:0]>15'b100010000000000))
                begin
                    addra4=6'b011010;
                    addrb4=6'b011011;
                end
            else if((x4[14:0]<=15'b100011000000000)&&(x4[14:0]>15'b100010100000000))
                begin
                    addra4=6'b011100;
                    addrb4=6'b011101;
                end
            else if((x4[14:0]<=15'b100011100000000)&&(x4[14:0]>15'b100011000000000))
                begin
                    addra4=6'b011110;
                    addrb4=6'b011111;
                end
            else if((x4[14:0]<=15'b100100000000000)&&(x4[14:0]>15'b100011100000000))
                begin
                    addra4=6'b100000;
                    addrb4=6'b100001;
                end
            else if((x4[14:0]<=15'b100100010000000)&&(x4[14:0]>15'b100100000000000))
                begin
                    addra4=6'b100010;
                    addrb4=6'b100011;
                end
            else if((x4[14:0]<=15'b100100100000000)&&(x4[14:0]>15'b100100010000000))
                begin
                    addra4=6'b100100;
                    addrb4=6'b100101;
                end
        end
        end
        always @(posedge aclk)
    begin
    if(x5[15:15]==1)
            begin
            if((x5[14:0]<=15'b100100010000000)&&(x5[14:0]>15'b100100000000000)) 
                begin
                    addra5=6'b000000;
                    addrb5=6'b000001;
                end
            else if((x5[14:0]<=15'b100100000000000)&&(x5[14:0]>15'b100011100000000))
                begin
                    addra5=6'b000010;
                    addrb5=6'b000011;
                end
            else if((x5[14:0]<=15'b100011100000000)&&(x5[14:0]>15'b100011000000000))
                begin
                    addra5=6'b000100;
                    addrb5=6'b000101;
                end
            else if((x5[14:0]<=15'b100011000000000)&&(x5[14:0]>15'b100010100000000))
                begin
                    addra5=6'b000110;
                    addrb5=6'b000111;
                end
            else if((x5[14:0]<=15'b100010100000000)&&(x5[14:0]>15'b100010000000000))
                begin
                    addra5=6'b001000;
                    addrb5=6'b001001;
                end
            else if((x5[14:0]<=15'b100010000000000)&&(x5[14:0]>15'b100001000000000))
                begin
                    addra5=6'b001010;
                    addrb5=6'b001011;
                end
            else if((x5[14:0]<=15'b100001000000000)&&(x5[14:0]>15'b100000000000000))
                begin
                    addra5=6'b001100;
                    addrb5=6'b001101;
                end
            else if((x5[14:0]<=15'b100000000000000)&&(x5[14:0]>15'b011110000000000))
                begin
                    addra5=6'b001110;
                    addrb5=6'b001111;
                end
            else if((x5[14:0]<=15'b011110000000000)&&(x5[14:0]>15'b000000000000000))
                begin
                    addra5=6'b010000;
                    addrb5=6'b010001;
                end
                end
    else
         begin
            if((x5[14:0]<=15'b011110000000000)&&(x5[14:0]>15'b000000000000000))
                begin
                    addra5=6'b010010;
                    addrb5=6'b010011;
                end
            else if((x5[14:0]<=15'b100000000000000)&&(x5>15'b011110000000000))
                begin
                    addra5=6'b010100;
                    addrb5=6'b010101;
                end
            else if((x5[14:0]<=15'b100001000000000)&&(x5>15'b100000000000000))
                begin
                    addra5=6'b010110;
                    addrb5=6'b010111;
                end
            else if((x5[14:0]<=15'b100010000000000)&&(x5[14:0]>15'b100001000000000))
                begin
                    addra5=6'b011000;
                    addrb5=6'b011001;
                end
            else if((x5[14:0]<=15'b100010100000000)&&(x5[14:0]>15'b100010000000000))
                begin
                    addra5=6'b011010;
                    addrb5=6'b011011;
                end
            else if((x5[14:0]<=15'b100011000000000)&&(x5[14:0]>15'b100010100000000))
                begin
                    addra5=6'b011100;
                    addrb5=6'b011101;
                end
            else if((x5[14:0]<=15'b100011100000000)&&(x5[14:0]>15'b100011000000000))
                begin
                    addra5=6'b011110;
                    addrb5=6'b011111;
                end
            else if((x5[14:0]<=15'b100100000000000)&&(x5[14:0]>15'b100011100000000))
                begin
                    addra5=6'b100000;
                    addrb5=6'b100001;
                end
            else if((x5[14:0]<=15'b100100010000000)&&(x5[14:0]>15'b100100000000000))
                begin
                    addra5=6'b100010;
                    addrb5=6'b100011;
                end
            else if((x5[14:0]<=15'b100100100000000)&&(x5[14:0]>15'b100100010000000))
                begin
                    addra5=6'b100100;
                    addrb5=6'b100101;
                end
        end
        end
        always @(posedge aclk)
    begin
    if(x6[15:15]==1)
            begin
            if((x6[14:0]<=15'b100100010000000)&&(x6[14:0]>15'b100100000000000)) 
                begin
                    addra6=6'b000000;
                    addrb6=6'b000001;
                end
            else if((x6[14:0]<=15'b100100000000000)&&(x6[14:0]>15'b100011100000000))
                begin
                    addra6=6'b000010;
                    addrb6=6'b000011;
                end
            else if((x6[14:0]<=15'b100011100000000)&&(x6[14:0]>15'b100011000000000))
                begin
                    addra6=6'b000100;
                    addrb6=6'b000101;
                end
            else if((x6[14:0]<=15'b100011000000000)&&(x6[14:0]>15'b100010100000000))
                begin
                    addra6=6'b000110;
                    addrb6=6'b000111;
                end
            else if((x6[14:0]<=15'b100010100000000)&&(x6[14:0]>15'b100010000000000))
                begin
                    addra6=6'b001000;
                    addrb6=6'b001001;
                end
            else if((x6[14:0]<=15'b100010000000000)&&(x6[14:0]>15'b100001000000000))
                begin
                    addra6=6'b001010;
                    addrb6=6'b001011;
                end
            else if((x6[14:0]<=15'b100001000000000)&&(x6[14:0]>15'b100000000000000))
                begin
                    addra6=6'b001100;
                    addrb6=6'b001101;
                end
            else if((x6[14:0]<=15'b100000000000000)&&(x6[14:0]>15'b011110000000000))
                begin
                    addra6=6'b001110;
                    addrb6=6'b001111;
                end
            else if((x6[14:0]<=15'b011110000000000)&&(x6[14:0]>15'b000000000000000))
                begin
                    addra6=6'b010000;
                    addrb6=6'b010001;
                end
                end
    else
         begin
            if((x6[14:0]<=15'b011110000000000)&&(x6[14:0]>15'b000000000000000))
                begin
                    addra6=6'b010010;
                    addrb6=6'b010011;
                end
            else if((x6[14:0]<=15'b100000000000000)&&(x6>15'b011110000000000))
                begin
                    addra6=6'b010100;
                    addrb6=6'b010101;
                end
            else if((x6[14:0]<=15'b100001000000000)&&(x6>15'b100000000000000))
                begin
                    addra6=6'b010110;
                    addrb6=6'b010111;
                end
            else if((x6[14:0]<=15'b100010000000000)&&(x6[14:0]>15'b100001000000000))
                begin
                    addra6=6'b011000;
                    addrb6=6'b011001;
                end
            else if((x6[14:0]<=15'b100010100000000)&&(x6[14:0]>15'b100010000000000))
                begin
                    addra6=6'b011010;
                    addrb6=6'b011011;
                end
            else if((x6[14:0]<=15'b100011000000000)&&(x6[14:0]>15'b100010100000000))
                begin
                    addra6=6'b011100;
                    addrb6=6'b011101;
                end
            else if((x6[14:0]<=15'b100011100000000)&&(x6[14:0]>15'b100011000000000))
                begin
                    addra6=6'b011110;
                    addrb6=6'b011111;
                end
            else if((x6[14:0]<=15'b100100000000000)&&(x6[14:0]>15'b100011100000000))
                begin
                    addra6=6'b100000;
                    addrb6=6'b100001;
                end
            else if((x6[14:0]<=15'b100100010000000)&&(x6[14:0]>15'b100100000000000))
                begin
                    addra6=6'b100010;
                    addrb6=6'b100011;
                end
            else if((x6[14:0]<=15'b100100100000000)&&(x6[14:0]>15'b100100010000000))
                begin
                    addra6=6'b100100;
                    addrb6=6'b100101;
                end
        end
        end
        always @(posedge aclk)
    begin
    if(x7[15:15]==1)
            begin
            if((x7[14:0]<=15'b100100010000000)&&(x7[14:0]>15'b100100000000000)) 
                begin
                    addra7=6'b000000;
                    addrb7=6'b000001;
                end
            else if((x7[14:0]<=15'b100100000000000)&&(x7[14:0]>15'b100011100000000))
                begin
                    addra7=6'b000010;
                    addrb7=6'b000011;
                end
            else if((x7[14:0]<=15'b100011100000000)&&(x7[14:0]>15'b100011000000000))
                begin
                    addra7=6'b000100;
                    addrb7=6'b000101;
                end
            else if((x7[14:0]<=15'b100011000000000)&&(x7[14:0]>15'b100010100000000))
                begin
                    addra7=6'b000110;
                    addrb7=6'b000111;
                end
            else if((x7[14:0]<=15'b100010100000000)&&(x7[14:0]>15'b100010000000000))
                begin
                    addra7=6'b001000;
                    addrb7=6'b001001;
                end
            else if((x7[14:0]<=15'b100010000000000)&&(x7[14:0]>15'b100001000000000))
                begin
                    addra7=6'b001010;
                    addrb7=6'b001011;
                end
            else if((x7[14:0]<=15'b100001000000000)&&(x7[14:0]>15'b100000000000000))
                begin
                    addra7=6'b001100;
                    addrb7=6'b001101;
                end
            else if((x7[14:0]<=15'b100000000000000)&&(x7[14:0]>15'b011110000000000))
                begin
                    addra7=6'b001110;
                    addrb7=6'b001111;
                end
            else if((x7[14:0]<=15'b011110000000000)&&(x7[14:0]>15'b000000000000000))
                begin
                    addra7=6'b010000;
                    addrb7=6'b010001;
                end
                end
    else
         begin
            if((x7[14:0]<=15'b011110000000000)&&(x7[14:0]>15'b000000000000000))
                begin
                    addra7=6'b010010;
                    addrb7=6'b010011;
                end
            else if((x7[14:0]<=15'b100000000000000)&&(x7>15'b011110000000000))
                begin
                    addra7=6'b010100;
                    addrb7=6'b010101;
                end
            else if((x7[14:0]<=15'b100001000000000)&&(x7>15'b100000000000000))
                begin
                    addra7=6'b010110;
                    addrb7=6'b010111;
                end
            else if((x7[14:0]<=15'b100010000000000)&&(x7[14:0]>15'b100001000000000))
                begin
                    addra7=6'b011000;
                    addrb7=6'b011001;
                end
            else if((x7[14:0]<=15'b100010100000000)&&(x7[14:0]>15'b100010000000000))
                begin
                    addra7=6'b011010;
                    addrb7=6'b011011;
                end
            else if((x7[14:0]<=15'b100011000000000)&&(x7[14:0]>15'b100010100000000))
                begin
                    addra7=6'b011100;
                    addrb7=6'b011101;
                end
            else if((x7[14:0]<=15'b100011100000000)&&(x7[14:0]>15'b100011000000000))
                begin
                    addra7=6'b011110;
                    addrb7=6'b011111;
                end
            else if((x7[14:0]<=15'b100100000000000)&&(x7[14:0]>15'b100011100000000))
                begin
                    addra7=6'b100000;
                    addrb7=6'b100001;
                end
            else if((x7[14:0]<=15'b100100010000000)&&(x7[14:0]>15'b100100000000000))
                begin
                    addra7=6'b100010;
                    addrb7=6'b100011;
                end
            else if((x7[14:0]<=15'b100100100000000)&&(x7[14:0]>15'b100100010000000))
                begin
                    addra7=6'b100100;
                    addrb7=6'b100101;
                end
        end
        end
    always @(posedge aclk)
    begin
    if(x8[15:15]==1)
            begin
            if((x8[14:0]<=15'b100100010000000)&&(x8[14:0]>15'b100100000000000)) 
                begin
                    addra8=6'b000000;
                    addrb8=6'b000001;
                end
            else if((x8[14:0]<=15'b100100000000000)&&(x8[14:0]>15'b100011100000000))
                begin
                    addra8=6'b000010;
                    addrb8=6'b000011;
                end
            else if((x8[14:0]<=15'b100011100000000)&&(x8[14:0]>15'b100011000000000))
                begin
                    addra8=6'b000100;
                    addrb8=6'b000101;
                end
            else if((x8[14:0]<=15'b100011000000000)&&(x8[14:0]>15'b100010100000000))
                begin
                    addra8=6'b000110;
                    addrb8=6'b000111;
                end
            else if((x8[14:0]<=15'b100010100000000)&&(x8[14:0]>15'b100010000000000))
                begin
                    addra8=6'b001000;
                    addrb8=6'b001001;
                end
            else if((x8[14:0]<=15'b100010000000000)&&(x8[14:0]>15'b100001000000000))
                begin
                    addra8=6'b001010;
                    addrb8=6'b001011;
                end
            else if((x8[14:0]<=15'b100001000000000)&&(x8[14:0]>15'b100000000000000))
                begin
                    addra8=6'b001100;
                    addrb8=6'b001101;
                end
            else if((x8[14:0]<=15'b100000000000000)&&(x8[14:0]>15'b011110000000000))
                begin
                    addra8=6'b001110;
                    addrb8=6'b001111;
                end
            else if((x8[14:0]<=15'b011110000000000)&&(x8[14:0]>15'b000000000000000))
                begin
                    addra8=6'b010000;
                    addrb8=6'b010001;
                end
                end
    else
         begin
            if((x8[14:0]<=15'b011110000000000)&&(x8[14:0]>15'b000000000000000))
                begin
                    addra8=6'b010010;
                    addrb8=6'b010011;
                end
            else if((x8[14:0]<=15'b100000000000000)&&(x8>15'b011110000000000))
                begin
                    addra8=6'b010100;
                    addrb8=6'b010101;
                end
            else if((x8[14:0]<=15'b100001000000000)&&(x8>15'b100000000000000))
                begin
                    addra8=6'b010110;
                    addrb8=6'b010111;
                end
            else if((x8[14:0]<=15'b100010000000000)&&(x8[14:0]>15'b100001000000000))
                begin
                    addra8=6'b011000;
                    addrb8=6'b011001;
                end
            else if((x8[14:0]<=15'b100010100000000)&&(x8[14:0]>15'b100010000000000))
                begin
                    addra8=6'b011010;
                    addrb8=6'b011011;
                end
            else if((x8[14:0]<=15'b100011000000000)&&(x8[14:0]>15'b100010100000000))
                begin
                    addra8=6'b011100;
                    addrb8=6'b011101;
                end
            else if((x8[14:0]<=15'b100011100000000)&&(x8[14:0]>15'b100011000000000))
                begin
                    addra8=6'b011110;
                    addrb8=6'b011111;
                end
            else if((x8[14:0]<=15'b100100000000000)&&(x8[14:0]>15'b100011100000000))
                begin
                    addra8=6'b100000;
                    addrb8=6'b100001;
                end
            else if((x8[14:0]<=15'b100100010000000)&&(x8[14:0]>15'b100100000000000))
                begin
                    addra8=6'b100010;
                    addrb8=6'b100011;
                end
            else if((x8[14:0]<=15'b100100100000000)&&(x8[14:0]>15'b100100010000000))
                begin
                    addra8=6'b100100;
                    addrb8=6'b100101;
                end
        end
        end
        always @(posedge aclk)
    begin
    if(x9[15:15]==1)
            begin
            if((x9[14:0]<=15'b100100010000000)&&(x9[14:0]>15'b100100000000000)) 
                begin
                    addra9=6'b000000;
                    addrb9=6'b000001;
                end
            else if((x9[14:0]<=15'b100100000000000)&&(x9[14:0]>15'b100011100000000))
                begin
                    addra9=6'b000010;
                    addrb9=6'b000011;
                end
            else if((x9[14:0]<=15'b100011100000000)&&(x9[14:0]>15'b100011000000000))
                begin
                    addra9=6'b000100;
                    addrb9=6'b000101;
                end
            else if((x9[14:0]<=15'b100011000000000)&&(x9[14:0]>15'b100010100000000))
                begin
                    addra9=6'b000110;
                    addrb9=6'b000111;
                end
            else if((x9[14:0]<=15'b100010100000000)&&(x9[14:0]>15'b100010000000000))
                begin
                    addra9=6'b001000;
                    addrb9=6'b001001;
                end
            else if((x9[14:0]<=15'b100010000000000)&&(x9[14:0]>15'b100001000000000))
                begin
                    addra9=6'b001010;
                    addrb9=6'b001011;
                end
            else if((x9[14:0]<=15'b100001000000000)&&(x9[14:0]>15'b100000000000000))
                begin
                    addra9=6'b001100;
                    addrb9=6'b001101;
                end
            else if((x9[14:0]<=15'b100000000000000)&&(x9[14:0]>15'b011110000000000))
                begin
                    addra9=6'b001110;
                    addrb9=6'b001111;
                end
            else if((x9[14:0]<=15'b011110000000000)&&(x9[14:0]>15'b000000000000000))
                begin
                    addra9=6'b010000;
                    addrb9=6'b010001;
                end
                end
    else
         begin
            if((x9[14:0]<=15'b011110000000000)&&(x9[14:0]>15'b000000000000000))
                begin
                    addra9=6'b010010;
                    addrb9=6'b010011;
                end
            else if((x9[14:0]<=15'b100000000000000)&&(x9>15'b011110000000000))
                begin
                    addra9=6'b010100;
                    addrb9=6'b010101;
                end
            else if((x9[14:0]<=15'b100001000000000)&&(x9>15'b100000000000000))
                begin
                    addra9=6'b010110;
                    addrb9=6'b010111;
                end
            else if((x9[14:0]<=15'b100010000000000)&&(x9[14:0]>15'b100001000000000))
                begin
                    addra9=6'b011000;
                    addrb9=6'b011001;
                end
            else if((x9[14:0]<=15'b100010100000000)&&(x9[14:0]>15'b100010000000000))
                begin
                    addra9=6'b011010;
                    addrb9=6'b011011;
                end
            else if((x9[14:0]<=15'b100011000000000)&&(x9[14:0]>15'b100010100000000))
                begin
                    addra9=6'b011100;
                    addrb9=6'b011101;
                end
            else if((x9[14:0]<=15'b100011100000000)&&(x9[14:0]>15'b100011000000000))
                begin
                    addra9=6'b011110;
                    addrb9=6'b011111;
                end
            else if((x9[14:0]<=15'b100100000000000)&&(x9[14:0]>15'b100011100000000))
                begin
                    addra9=6'b100000;
                    addrb9=6'b100001;
                end
            else if((x9[14:0]<=15'b100100010000000)&&(x9[14:0]>15'b100100000000000))
                begin
                    addra9=6'b100010;
                    addrb9=6'b100011;
                end
            else if((x9[14:0]<=15'b100100100000000)&&(x9[14:0]>15'b100100010000000))
                begin
                    addra9=6'b100100;
                    addrb9=6'b100101;
                end
        end
        end  
endmodule
